* DC model fitted to graphs in datasheet

.SUBCKT aptf1616lseezgkqbkc-dc A R G B
D1 A R red
D2 A G green
D3 A B blue

.MODEL red D
+ IS=8.005438771378796e-11
+ N=3.9378148558540444
+ RS=1.7463723493295458
+ TNOM=295

.MODEL green D
+ IS=7.856521889175404e-11
+ N=6.06505638107386
+ RS=8.94568304574287
+ TNOM=295

.MODEL blue D
+ IS=8.880842070259583e-11
+ N=6.000925797457152
+ RS=12.976314392284344
+ TNOM=295

.ENDS
